`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BcTuTm10kQEWxearr2PjwSnO7Ywl9LEsP58yPequqaNPFEVPpVJ9gd6Vp8XC+Gno
1iaKyvw/NnrnWTZ+o61arRr93F6xAiZuvAWb2kcTPY0sBM8FqkulToTh8mU18nWH
gHtP5D4qAGe4WA1uhy/zjQ==
`protect END_PROTECTED
