library verilog;
use verilog.vl_types.all;
entity float_pack_tb is
end float_pack_tb;
