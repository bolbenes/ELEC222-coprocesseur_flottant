package float_pack; 
// Ajouter ici les définition des fonctions
   // utilisée par votre coprocesseur
   parameter Nm =`TB_MANT_SIZE;
   parameter Ne = `TB_EXP_SIZE;
   `include "../find_first_bit_one.sv"
   typedef struct packed 
		  {
		     logic signe;
		     logic [Ne-1:0] exponent;
		     logic [Nm-1:0] mantisse;
		  } float;
   
   typedef struct packed 
		  {
		     logic signe;
		     logic [8-1:0] exponent;
		     logic [23-1:0]  mantisse;
		  } float_ieee;

   function float_ieee real2float_ieee ( input shortreal real_in);
	 return ($shortrealtobits(real_in));
   endfunction // real2float_ieee
   
   function shortreal float_ieee2real ( input float_ieee float_in);
      return ($bitstoshortreal(float_in));
   endfunction // float_ieee2real

   function float real2float (input shortreal real_in);
	return (float_ieee2float($shortrealtobits(real_in)));
   endfunction // real2float

   function shortreal float2real (input float float_in);
     return $bitstoshortreal(float2float_ieee(float_in));
   endfunction // float2real
   

   // condition: float: moins de bits que float_ieee
   function float_ieee float2float_ieee(input float float_in);
      
      float_ieee result;
      
     begin
	result.exponent = float_in.exponent+127-(2**(Ne-1)-1);
	result.mantisse = '0;
	result.mantisse[22:22-(Nm-1)] = float_in.mantisse;
	result.signe = float_in.signe;
	return result;
     end
   endfunction // float2float_ieee
   
   function float float_ieee2float(input float_ieee float_in);
      
      integer exposant;
      float result;
      
      begin
	 exposant = float_in.exponent - 127;
	 if(exposant <= 2**(Ne-1)-1 && exposant >= -2**(Ne-1)+2)
	   begin
	      result.exponent = exposant + 2**(Ne-1)-1;
	      result.mantisse = float_in.mantisse[22:22-(Nm-1)];
	   end
	 else if(exposant > 2**(Ne-1)-1)
	   begin
	      result.exponent = 2**Ne-2;
	      result.mantisse = '1;
	   end
	 else if(exposant < -2**(Ne-1)+2)
	   begin
	      result.exponent = '0;
	      result.mantisse = '0;
	   end
	 result.signe = float_in.signe;
	 return result;
      end
   endfunction // float_ieee2float
   
   function float float_mul(input float A, input float B);
      
      float result,max_exposant,min_exposant;
      logic [Nm:0] mantisse_max, mantisse_min;
      logic [2*Nm:0] mantisse_result;
            
      begin
	 // on calcule le signe
	 result.signe = A.signe + B.signe;
	 // on calcule l'exposant
	 result.exponent = A.exponent + B.exponent + (2**(Ne-1)-1);
	 //calcul de la mantisse
	 if (A.exponent < B.exponent)
	   begin
	      mantisse_max = {1,B.mantisse};
	      mantisse_min ={1,A.mantisse};
	      mantisse_result = mantisse_max * (mantisse_min >> (A.exponent - B.exponent));// on décale la mantisse de l'écart entre les exposants
	   end
	 else
	   begin
	      mantisse_max = {1,A.mantisse};
	      mantisse_min ={1,B.mantisse};
	      mantisse_result = mantisse_max * (mantisse_min >> (A.exponent - B.exponent));// on décale la mantisse de l'écart entre les exposants
	   end // else: !if(A.exponent < B.exponent)
	 if (mantisse_result*2**(-2*Nm)>=2)
	   begin
	      result.exponent = result.exponent +1;
	      result.mantisse = (mantisse_result[2*Nm-1:Nm-1]>>1);
	   end
	 else
	   result.mantisse = mantisse_result[2*Nm-1:Nm-1];
	 
	 return result; 
      end
   endfunction
   
   logic[23:0] findfirst1;
   logic [4:0] resultfirst1;
	
   function float float_add(input float A, input float B);
      return float_add_sub(A,B,0);
   endfunction
   
   function float float_add_sub(input float A, input float B, logic add_sub); // add: add_sub=0, sub: add_sub=1
      logic [7:0] exp_difference;
      logic [24:-2] shifted_mantisse;
      logic [24:-2] temp1, temp2; // les mantisses qu'on additionne
      logic [25:-2] result_mantisse_unnorm;
      logic [23:0] mantisse_to_check;
      logic [4:0] result_first_one; 
      logic [47:-2] temp_shift;
      logic [47:0] temp_mantisse;
      logic [9:0]  result_exponent;
      logic [22:0] result_mantisse;
      logic 	   result_signe;
      float Aa,Bb;
      
      logic 	   subtrahend = 0; // 0 signifie, que B est le subtrahend, 1 signifie que A est le subtrahend
      begin
	 //$display("A.sign = %b\nA.mantisse = %b\nA.exponent = %b\n",A.signe,A.mantisse,A.exponent);
	 //$display("B.sign = %b\nB.mantisse = %b\nB.exponent = %b\n",B.signe,B.mantisse,B.exponent);
	 
	 if({A.exponent,A.mantisse} <= {B.exponent,B.mantisse})
	   begin
	      Aa = B;
	      Bb = A;
	   subtrahend = 1;
	   end
	 else
	   begin
	      Aa = A;
	      Bb = B;
	   end // else: !if(A.exponent <= B.exponent)

	 if({Bb.mantisse,Bb.exponent} == '0)
	   return Aa;
	 
	 
	 //$display("\nNouveau calcul\nAa.signe %b\nAa.mantisse %b\nAa.exponent %b\nBb.signe %b\nBb.mantisse %b\nBb.exponent %b",Aa.signe,Aa.mantisse,Aa.exponent,Bb.signe,Bb.mantisse,Bb.exponent);
	 
	 exp_difference = Aa.exponent-Bb.exponent;
	 if(exp_difference > Nm-1)
	   return Aa;
         temp_shift = '0;
         temp_shift[23] = 1;
         temp_shift[22:0]= Bb.mantisse;

	 //$display("\nexp_difference: %b",exp_difference);
	 shifted_mantisse = '0;
         shifted_mantisse[23:-2] = temp_shift[23+exp_difference-:26];
	 //$display("Aa.mantisse:\t\t\t %b",Aa.mantisse);
	 //$display("shifted mantisse de Bb:\t %b",shifted_mantisse);
	 temp1 = {2'b01, Aa.mantisse,2'b0};
	 //$display("mantisse de Aa:\t\t %b\n",temp1);
	 temp2 = shifted_mantisse;
	 
	 
	 if(add_sub == 0) // add
	   begin
	      result_signe = Aa.signe;
	      if(Aa.signe == Bb.signe)
		begin
		   result_mantisse_unnorm = temp1+temp2;
		end
	      else
		begin
		   result_mantisse_unnorm = temp1-temp2;
		end
	   end // if (add_sub == 0)
	 else // sub
	   begin
	      if(Aa.signe == 0)
		begin
		   result_signe = subtrahend;		   
		end
	      else
		begin
		   result_signe = ~subtrahend;
		end
	      if(Aa.signe == Bb.signe)
		begin
		   result_mantisse_unnorm = temp1-temp2;
		end
	      else
		begin
		   result_mantisse_unnorm = temp1+temp2;
		end	      
	   end // else: !if(add_sub == 0)

	 //$display("result_mantisse_unnorm: \t%b",result_mantisse_unnorm);
	 //$display("result_signe: %b",result_signe);
	 
    
	 resultfirst1 = find_first_bit_one(result_mantisse_unnorm[25:2]);
         //$display("first 1: %d",resultfirst1);

	 if(resultfirst1 == 5'b0 && result_mantisse_unnorm[2:0] == 3'b0)
	   begin
	      result_mantisse = '0;
	      Aa.exponent = '0;
	   end
	 else
	   begin
	      result_mantisse_unnorm = result_mantisse_unnorm << (25-resultfirst1-1);
	      result_mantisse = result_mantisse_unnorm[25-:23];
	      result_exponent = Aa.exponent - (21-resultfirst1);
	      if(result_exponent[9] == 1 || result_exponent == '0)
		begin
		   result_exponent = '0;
		   result_mantisse = '0;
		end
	      else if(result_exponent[8:0] > 2**(Ne)-2)
		begin
		   result_exponent = '1;
		   result_mantisse = '0;
		end
	   
	      Aa.exponent = result_exponent;
	   end
	 /*
         temp_mantisse = '0;
         temp_mantisse[47:24]=result_mantisse;
         result_mantisse = '0;
	 	 
         result_mantisse = temp_mantisse[(47-(24-resultfirst1))-:24];
	 */
	 //$display("result_mantisse = %b", result_mantisse);
	 
         
         Aa.signe = result_signe;
         Aa.mantisse = result_mantisse;
	 //$display("Aa.sign = %b\nAa.mantisse = %b\nAa.exponent = %b\n",Aa.signe,Aa.mantisse,Aa.exponent);

         return Aa;
      end
   endfunction // float_add_sub
endpackage : float_pack
   
   